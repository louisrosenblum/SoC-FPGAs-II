ROM_1_PORT_inst : ROM_1_PORT PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
